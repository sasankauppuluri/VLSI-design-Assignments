magic
tech scmos
timestamp 1613748099
<< nwell >>
rect -13 -7 15 30
<< ntransistor >>
rect 0 -26 2 -16
<< ptransistor >>
rect 0 -1 2 24
<< ndiffusion >>
rect -1 -26 0 -16
rect 2 -26 3 -16
<< pdiffusion >>
rect -1 -1 0 24
rect 2 -1 3 24
<< ndcontact >>
rect -6 -26 -1 -16
rect 3 -26 8 -16
<< pdcontact >>
rect -6 -1 -1 24
rect 3 -1 8 24
<< polysilicon >>
rect 0 24 2 27
rect 0 -16 2 -1
rect 0 -30 2 -26
<< polycontact >>
rect -6 -13 0 -8
<< metal1 >>
rect -13 29 15 35
rect -6 24 -1 29
rect 3 -8 8 -1
rect -18 -13 -6 -8
rect 3 -13 21 -8
rect 3 -16 8 -13
rect -6 -32 -1 -26
rect -13 -36 15 -32
<< labels >>
rlabel metal1 -13 29 15 35 5 vdd
rlabel metal1 -13 -36 15 -32 1 gnd
rlabel metal1 -18 -13 0 -8 1 input
rlabel metal1 3 -13 21 -8 1 output
<< end >>
