magic
tech scmos
timestamp 1613661510
<< metal1 >>
rect 5 104 75 112
rect 6 0 75 4
use cmosinverter1  cmosinverter1_0
timestamp 1613660981
transform 1 0 8 0 1 42
box -8 -42 33 70
use cmosinverter1  cmosinverter1_1
timestamp 1613660981
transform 1 0 49 0 1 42
box -8 -42 33 70
<< labels >>
rlabel metal1 5 104 75 112 5 vdd
rlabel metal1 6 0 75 4 1 gnd
rlabel space 0 33 19 38 1 input
rlabel space 68 33 82 38 1 output
<< end >>
