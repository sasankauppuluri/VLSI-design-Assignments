magic
tech scmos
timestamp 1613758697
<< metal1 >>
rect -7 -19 2 28
rect -7 -24 39 -19
rect 624 -24 634 28
use inverter5  inverter5_0
array 0 15 39 0 0 71
timestamp 1613748099
transform 1 0 18 0 1 36
box -18 -36 21 35
use inverter5  inverter5_1
array 0 14 -39 0 0 -71
timestamp 1613748099
transform -1 0 60 0 -1 -32
box -18 -36 21 35
<< end >>
