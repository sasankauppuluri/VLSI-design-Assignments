magic
tech scmos
timestamp 1613749228
<< metal1 >>
rect -17 -55 -12 25
rect 612 20 623 25
rect 618 -55 623 20
rect -17 -60 27 -55
rect 612 -60 623 -55
use inverter5  inverter5_0
array 0 15 39 0 0 71
timestamp 1613748099
transform 1 0 6 0 1 33
box -18 -36 21 35
use inverter5  inverter5_1
array 0 14 -39 0 0 71
timestamp 1613748099
transform -1 0 48 0 1 -47
box -18 -36 21 35
<< end >>
